module bitwiseand(out,x,y);
    input [31:0] x;
    input [31:0] y;
    output [31:0] out;

    and b0(out[0], x[0], y[0]);
    and b1(out[1], x[1], y[1]);
    and b2(out[2], x[2], y[2]);
    and b3(out[3], x[3], y[3]);
    and b4(out[4], x[4], y[4]);
    and b5(out[5], x[5], y[5]);
    and b6(out[6], x[6], y[6]);
    and b7(out[7], x[7], y[7]);
    and b8(out[8], x[8], y[8]);
    and b9(out[9], x[9], y[9]);
    and b10(out[10], x[10], y[10]);
    and b11(out[11], x[11], y[11]);
    and b12(out[12], x[12], y[12]);
    and b13(out[13], x[13], y[13]);
    and b14(out[14], x[14], y[14]);
    and b15(out[15], x[15], y[15]);
    and b16(out[16], x[16], y[16]);
    and b17(out[17], x[17], y[17]);
    and b18(out[18], x[18], y[18]);
    and b19(out[19], x[19], y[19]);
    and b20(out[20], x[20], y[20]);
    and b21(out[21], x[21], y[21]);
    and b22(out[22], x[22], y[22]);
    and b23(out[23], x[23], y[23]);
    and b24(out[24], x[24], y[24]);
    and b25(out[25], x[25], y[25]);
    and b26(out[26], x[26], y[26]);
    and b27(out[27], x[27], y[27]);
    and b28(out[28], x[28], y[28]);
    and b29(out[29], x[29], y[29]);
    and b30(out[30], x[30], y[30]);
    and b31(out[31], x[31], y[31]);
endmodule

module bitwiseor(out,x,y);
    input [31:0] x;
    input [31:0] y;
    output [31:0] out;

    or b0(out[0], x[0], y[0]);
    or b1(out[1], x[1], y[1]);
    or b2(out[2], x[2], y[2]);
    or b3(out[3], x[3], y[3]);
    or b4(out[4], x[4], y[4]);
    or b5(out[5], x[5], y[5]);
    or b6(out[6], x[6], y[6]);
    or b7(out[7], x[7], y[7]);
    or b8(out[8], x[8], y[8]);
    or b9(out[9], x[9], y[9]);
    or b10(out[10], x[10], y[10]);
    or b11(out[11], x[11], y[11]);
    or b12(out[12], x[12], y[12]);
    or b13(out[13], x[13], y[13]);
    or b14(out[14], x[14], y[14]);
    or b15(out[15], x[15], y[15]);
    or b16(out[16], x[16], y[16]);
    or b17(out[17], x[17], y[17]);
    or b18(out[18], x[18], y[18]);
    or b19(out[19], x[19], y[19]);
    or b20(out[20], x[20], y[20]);
    or b21(out[21], x[21], y[21]);
    or b22(out[22], x[22], y[22]);
    or b23(out[23], x[23], y[23]);
    or b24(out[24], x[24], y[24]);
    or b25(out[25], x[25], y[25]);
    or b26(out[26], x[26], y[26]);
    or b27(out[27], x[27], y[27]);
    or b28(out[28], x[28], y[28]);
    or b29(out[29], x[29], y[29]);
    or b30(out[30], x[30], y[30]);
    or b31(out[31], x[31], y[31]);
endmodule

module bitwisenot(out, x);
    input [31:0] x; // 32-bit input
    output [31:0] out; // 32-bit output

    not n0(out[0], x[0]);
    not n1(out[1], x[1]);
    not n2(out[2], x[2]);
    not n3(out[3], x[3]);
    not n4(out[4], x[4]);
    not n5(out[5], x[5]);
    not n6(out[6], x[6]);
    not n7(out[7], x[7]);
    not n8(out[8], x[8]);
    not n9(out[9], x[9]);
    not n10(out[10], x[10]);
    not n11(out[11], x[11]);
    not n12(out[12], x[12]);
    not n13(out[13], x[13]);
    not n14(out[14], x[14]);
    not n15(out[15], x[15]);
    not n16(out[16], x[16]);
    not n17(out[17], x[17]);
    not n18(out[18], x[18]);
    not n19(out[19], x[19]);
    not n20(out[20], x[20]);
    not n21(out[21], x[21]);
    not n22(out[22], x[22]);
    not n23(out[23], x[23]);
    not n24(out[24], x[24]);
    not n25(out[25], x[25]);
    not n26(out[26], x[26]);
    not n27(out[27], x[27]);
    not n28(out[28], x[28]);
    not n29(out[29], x[29]);
    not n30(out[30], x[30]);
    not n31(out[31], x[31]);
endmodule
